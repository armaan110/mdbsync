library verilog;
use verilog.vl_types.all;
entity MDP3_Parser_tb is
end MDP3_Parser_tb;
